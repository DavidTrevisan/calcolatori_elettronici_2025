library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package lfsr_pkg is
	function lfsr(x : in std_logic_vector) return std_logic_vector;
end lfsr_pkg;

library ieee;
use ieee.std_logic_1164.all;

package body lfsr_pkg is
	function get_poly(n : in integer) return std_logic_vector;

	function lfsr_int(x : in std_logic_vector) return std_logic_vector is
		variable poly		: std_logic_vector(63 downto 0);
		variable res		: std_logic_vector(x'range);
	begin
		if x'length < 1 or x'length > 64 then
			return x;
		elsif x'length < 2 then
			return not x;
		elsif x(x'right) = '1' then
			poly := get_poly(x'length);
			res := ('0' & x(x'left downto x'right + 1)) xor poly(x'length - 1 downto 0);
		else
			res := ('0' & x(x'left downto x'right + 1));
		end if;
		return res;
	end function lfsr_int;

	function lfsr(x : in std_logic_vector) return std_logic_vector is
	begin
		if x'length <= 64 then
			return lfsr_int(x);
		elsif x'length <= (64 + 63) then
			return lfsr_int(x(x'left downto 64)) & lfsr_int(x(63 downto 0));
		elsif x'length <= (64 + 63 + 62) then
			return
				lfsr_int(x(x'left downto 64 + 63)) &
				lfsr_int(x(64 + 63 - 1 downto 64)) &
				lfsr_int(x(63 downto 0));
		elsif x'length <= (64 + 63 + 62 + 61) then
			return
				lfsr_int(x(x'left downto 64 + 63 + 62)) &
				lfsr_int(x(64 + 63 + 62 - 1 downto 64 + 63)) &
				lfsr_int(x(64 + 63 - 1 downto 64)) &
				lfsr_int(x(63 downto 0));
		else
			return x;
		end if;
	end function lfsr;

	function get_poly(n : in integer) return std_logic_vector is
		type array_of_slv is array (natural range <>) of std_logic_vector(63 downto 0);
		constant polys		: array_of_slv := (
			"XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",	-- 0 invalid
			"XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",	-- 1 invalid
			"0000000000000000000000000000000000000000000000000000000000000011",	-- 2
			"0000000000000000000000000000000000000000000000000000000000000101",	-- 3
			"0000000000000000000000000000000000000000000000000000000000001001",	-- 4
			"0000000000000000000000000000000000000000000000000000000000010010",	-- 5
			"0000000000000000000000000000000000000000000000000000000000100001",	-- 6
			"0000000000000000000000000000000000000000000000000000000001000001",	-- 7
			"0000000000000000000000000000000000000000000000000000000010001110",	-- 8
			"0000000000000000000000000000000000000000000000000000000100001000",	-- 9
			"0000000000000000000000000000000000000000000000000000001000000100",	-- 10
			"0000000000000000000000000000000000000000000000000000010000000010",	-- 11
			"0000000000000000000000000000000000000000000000000000100000101001",	-- 12
			"0000000000000000000000000000000000000000000000000001000000001101",	-- 13
			"0000000000000000000000000000000000000000000000000010000000010101",	-- 14
			"0000000000000000000000000000000000000000000000000100000000000001",	-- 15
			"0000000000000000000000000000000000000000000000001000000000010110",	-- 16
			"0000000000000000000000000000000000000000000000010000000000000100",	-- 17
			"0000000000000000000000000000000000000000000000100000000000010011",	-- 18
			"0000000000000000000000000000000000000000000001000000000000010011",	-- 19
			"0000000000000000000000000000000000000000000010000000000000000100",	-- 20
			"0000000000000000000000000000000000000000000100000000000000000010",	-- 21
			"0000000000000000000000000000000000000000001000000000000000000001",	-- 22
			"0000000000000000000000000000000000000000010000000000000000010000",	-- 23
			"0000000000000000000000000000000000000000100000000000000000001101",	-- 24
			"0000000000000000000000000000000000000001000000000000000000000100",	-- 25
			"0000000000000000000000000000000000000010000000000000000000100011",	-- 26
			"0000000000000000000000000000000000000100000000000000000000010011",	-- 27
			"0000000000000000000000000000000000001000000000000000000000000100",	-- 28
			"0000000000000000000000000000000000010000000000000000000000000010",	-- 29
			"0000000000000000000000000000000000100000000000000000000000101001",	-- 30
			"0000000000000000000000000000000001000000000000000000000000000100",	-- 31
			"0000000000000000000000000000000010000000000000000000000001010111",	-- 32
			"0000000000000000000000000000000100000000000000000000000000101001",	-- 33
			"0000000000000000000000000000001000000000000000000000000001110011",	-- 34
			"0000000000000000000000000000010000000000000000000000000000000010",	-- 35
			"0000000000000000000000000000100000000000000000000000000000111011",	-- 36
			"0000000000000000000000000001000000000000000000000000000000011111",	-- 37
			"0000000000000000000000000010000000000000000000000000000000110001",	-- 38
			"0000000000000000000000000100000000000000000000000000000000001000",	-- 39
			"0000000000000000000000001000000000000000000000000000000000011100",	-- 40
			"0000000000000000000000010000000000000000000000000000000000000100",	-- 41
			"0000000000000000000000100000000000000000000000000000000000011111",	-- 42
			"0000000000000000000001000000000000000000000000000000000000101100",	-- 43
			"0000000000000000000010000000000000000000000000000000000000110010",	-- 44
			"0000000000000000000100000000000000000000000000000000000000001101",	-- 45
			"0000000000000000001000000000000000000000000000000000000010010111",	-- 46
			"0000000000000000010000000000000000000000000000000000000000010000",	-- 47
			"0000000000000000100000000000000000000000000000000000000001011011",	-- 48
			"0000000000000001000000000000000000000000000000000000000000111000",	-- 49
			"0000000000000010000000000000000000000000000000000000000000001110",	-- 50
			"0000000000000100000000000000000000000000000000000000000000100101",	-- 51
			"0000000000001000000000000000000000000000000000000000000000000100",	-- 52
			"0000000000010000000000000000000000000000000000000000000000100011",	-- 53
			"0000000000100000000000000000000000000000000000000000000000111110",	-- 54
			"0000000001000000000000000000000000000000000000000000000000100011",	-- 55
			"0000000010000000000000000000000000000000000000000000000001001010",	-- 56
			"0000000100000000000000000000000000000000000000000000000000010110",	-- 57
			"0000001000000000000000000000000000000000000000000000000000110001",	-- 58
			"0000010000000000000000000000000000000000000000000000000000111101",	-- 59
			"0000100000000000000000000000000000000000000000000000000000000001",	-- 60
			"0001000000000000000000000000000000000000000000000000000000010011",	-- 61
			"0010000000000000000000000000000000000000000000000000000000110100",	-- 62
			"0100000000000000000000000000000000000000000000000000000000000001",	-- 63
			"1000000000000000000000000000000000000000000000000000000000001101"	-- 64
		);

		variable idx		: natural;
		variable poly		: std_logic_vector(n - 1 downto 0);

	begin
		return polys(n);
	end function get_poly;
end lfsr_pkg;

